magic
tech sky130A
magscale 1 2
timestamp 1741188478
<< nwell >>
rect -696 -1219 696 1219
<< pmos >>
rect -500 -1000 500 1000
<< pdiff >>
rect -558 988 -500 1000
rect -558 -988 -546 988
rect -512 -988 -500 988
rect -558 -1000 -500 -988
rect 500 988 558 1000
rect 500 -988 512 988
rect 546 -988 558 988
rect 500 -1000 558 -988
<< pdiffc >>
rect -546 -988 -512 988
rect 512 -988 546 988
<< nsubdiff >>
rect -660 1149 -564 1183
rect 564 1149 660 1183
rect -660 1087 -626 1149
rect 626 1087 660 1149
rect -660 -1149 -626 -1087
rect 626 -1149 660 -1087
rect -660 -1183 -564 -1149
rect 564 -1183 660 -1149
<< nsubdiffcont >>
rect -564 1149 564 1183
rect -660 -1087 -626 1087
rect 626 -1087 660 1087
rect -564 -1183 564 -1149
<< poly >>
rect -500 1081 500 1097
rect -500 1047 -484 1081
rect 484 1047 500 1081
rect -500 1000 500 1047
rect -500 -1047 500 -1000
rect -500 -1081 -484 -1047
rect 484 -1081 500 -1047
rect -500 -1097 500 -1081
<< polycont >>
rect -484 1047 484 1081
rect -484 -1081 484 -1047
<< locali >>
rect -660 1149 -564 1183
rect 564 1149 660 1183
rect -660 1087 -626 1149
rect 626 1087 660 1149
rect -500 1047 -484 1081
rect 484 1047 500 1081
rect -546 988 -512 1004
rect -546 -1004 -512 -988
rect 512 988 546 1004
rect 512 -1004 546 -988
rect -500 -1081 -484 -1047
rect 484 -1081 500 -1047
rect -660 -1149 -626 -1087
rect 626 -1149 660 -1087
rect -660 -1183 -564 -1149
rect 564 -1183 660 -1149
<< viali >>
rect -484 1047 484 1081
rect -546 -988 -512 988
rect 512 -988 546 988
rect -484 -1081 484 -1047
<< metal1 >>
rect -496 1081 496 1087
rect -496 1047 -484 1081
rect 484 1047 496 1081
rect -496 1041 496 1047
rect -552 988 -506 1000
rect -552 -988 -546 988
rect -512 -988 -506 988
rect -552 -1000 -506 -988
rect 506 988 552 1000
rect 506 -988 512 988
rect 546 -988 552 988
rect 506 -1000 552 -988
rect -496 -1047 496 -1041
rect -496 -1081 -484 -1047
rect 484 -1081 496 -1047
rect -496 -1087 496 -1081
<< properties >>
string FIXED_BBOX -643 -1166 643 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
