* NGSPICE file created from OFC_parax.ext - technology: sky130A

.subckt OFC_parax VDD GND IN+ IN- OUT
X0 VDD.t8 Vp.t1 GND.t11 sky130_fd_pr__res_xhigh_po_0p35 l=5
X1 VDD.t3 G.t2 D10.t2 VDD.t2 sky130_fd_pr__pfet_01v8 ad=7.395 pd=51.58 as=7.395 ps=51.58 w=25.5 l=1
X2 w_1686_7818.t20 IN+.t0 D1.t3 w_1686_7818.t19 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X3 VDD.t1 Vp.t2 a_3651_12640# VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=5
X4 Vc.t0 GND.t5 GND.t4 sky130_fd_pr__res_xhigh_po_0p35 l=3.15
X5 w_1686_7818.t2 IN-.t0 D2.t4 w_1686_7818.t1 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X6 w_1686_7818.t4 IN-.t1 D2.t3 w_1686_7818.t3 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X7 Vp.t0 GND.t1 GND.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1.86
X8 VDD.t7 Vc.t1 GND.t10 sky130_fd_pr__res_xhigh_po_0p35 l=5
X9 D2.t6 Vc.t2 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=10
X10 VDD.t6 G.t3 D9.t2 VDD.t5 sky130_fd_pr__pfet_01v8 ad=7.395 pd=51.58 as=7.395 ps=51.58 w=25.5 l=1
X11 w_1686_7818.t18 IN+.t1 D1.t2 w_1686_7818.t17 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X12 w_1686_7818.t6 IN-.t2 D2.t2 w_1686_7818.t5 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X13 D10.t1 Vc.t3 OUT.t1 D10.t0 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=5
X14 w_1686_7818.t16 IN+.t2 D1.t4 w_1686_7818.t15 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X15 a_3651_12640# Vp.t3 w_1686_7818.t0 VDD.t4 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=5
X16 D9.t1 Vc.t4 G.t0 D9.t0 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=5
X17 w_1686_7818.t14 IN+.t3 D1.t5 w_1686_7818.t13 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X18 w_1686_7818.t8 IN-.t3 D2.t1 w_1686_7818.t7 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X19 G.t1 Vc.t5 D1.t1 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=2
X20 OUT.t0 Vc.t6 D2.t5 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=2
X21 w_1686_7818.t10 IN-.t4 D2.t0 w_1686_7818.t9 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X22 w_1686_7818.t12 IN+.t4 D1.t6 w_1686_7818.t11 sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X23 D1.t0 Vc.t7 GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=10
R0 VDD.n19 VDD.n13 10383.5
R1 VDD.n16 VDD.n14 10383.5
R2 VDD.n8 VDD.n2 10383.5
R3 VDD.n6 VDD.n5 10383.5
R4 VDD.n31 VDD.n29 4560
R5 VDD.n34 VDD.n33 4560
R6 VDD.n42 VDD.n40 4560
R7 VDD.n45 VDD.n44 4560
R8 VDD.n17 VDD.n13 3087.69
R9 VDD.n18 VDD.n14 3087.69
R10 VDD.n5 VDD.n4 3087.69
R11 VDD.n8 VDD.n7 3087.69
R12 VDD.n20 VDD.n12 1107.58
R13 VDD.n15 VDD.n12 1107.58
R14 VDD.n15 VDD.n11 1107.58
R15 VDD.n9 VDD.n1 1107.58
R16 VDD.n3 VDD.n1 1107.58
R17 VDD.n3 VDD.n0 1107.58
R18 VDD.n10 VDD.n0 902.898
R19 VDD.n21 VDD.n20 748.705
R20 VDD.n30 VDD.n26 486.401
R21 VDD.n30 VDD.n27 486.401
R22 VDD.n41 VDD.n37 486.401
R23 VDD.n41 VDD.n38 486.401
R24 VDD.n46 VDD.n38 460.425
R25 VDD.n35 VDD.n27 459.125
R26 VDD.n36 VDD.n26 441.337
R27 VDD.n47 VDD.n37 439.079
R28 VDD.n32 VDD.n31 421.394
R29 VDD.n34 VDD.n28 421.394
R30 VDD.n43 VDD.n42 421.394
R31 VDD.n45 VDD.n39 421.394
R32 VDD.n21 VDD.n11 294.68
R33 VDD.n10 VDD.n9 174.804
R34 VDD.n50 VDD.t1 48.1635
R35 VDD.n22 VDD.t7 43.7072
R36 VDD.n51 VDD.t8 42.6337
R37 VDD.n13 VDD.n12 37.0005
R38 VDD.n14 VDD.n11 37.0005
R39 VDD.n9 VDD.n8 37.0005
R40 VDD.n5 VDD.n3 37.0005
R41 VDD.n29 VDD.n26 10.8829
R42 VDD.n31 VDD.n30 10.8829
R43 VDD.n33 VDD.n27 10.8829
R44 VDD.n35 VDD.n34 10.8829
R45 VDD.n40 VDD.n37 10.8829
R46 VDD.n42 VDD.n41 10.8829
R47 VDD.n44 VDD.n38 10.8829
R48 VDD.n46 VDD.n45 10.8829
R49 VDD.n29 VDD.n28 9.85419
R50 VDD.n33 VDD.n32 9.85419
R51 VDD.n40 VDD.n39 9.85419
R52 VDD.n44 VDD.n43 9.85419
R53 VDD.n24 VDD.t6 9.05168
R54 VDD.n23 VDD.t3 9.05168
R55 VDD.n47 VDD.n46 5.7605
R56 VDD.n36 VDD.n35 4.8005
R57 VDD.n25 VDD.n10 3.1911
R58 VDD.n48 VDD.n36 2.79929
R59 VDD.n48 VDD.n47 2.4723
R60 VDD.n22 VDD.n21 2.40429
R61 VDD.n20 VDD.n19 2.37229
R62 VDD.n16 VDD.n15 2.37229
R63 VDD.n6 VDD.n1 2.37229
R64 VDD.n2 VDD.n0 2.37229
R65 VDD.n19 VDD.n18 1.66713
R66 VDD.n17 VDD.n16 1.66713
R67 VDD.n4 VDD.n2 1.66713
R68 VDD.n7 VDD.n6 1.66713
R69 VDD.n51 VDD.n50 1.40748
R70 VDD.n24 VDD.n23 1.39943
R71 VDD.n50 VDD.n49 1.01822
R72 VDD.t4 VDD.n28 1.00665
R73 VDD.n32 VDD.t4 1.00665
R74 VDD.t0 VDD.n39 1.00665
R75 VDD.n43 VDD.t0 1.00665
R76 VDD.n18 VDD.t2 0.706287
R77 VDD.t2 VDD.n17 0.706287
R78 VDD.n7 VDD.t5 0.706287
R79 VDD.n4 VDD.t5 0.706287
R80 VDD.n25 VDD.n24 0.530238
R81 VDD.n23 VDD.n22 0.419511
R82 VDD VDD.n51 0.332397
R83 VDD.n49 VDD.n48 0.201265
R84 VDD.n49 VDD.n25 0.153517
R85 Vp.n1 Vp.t1 43.2783
R86 Vp.n1 Vp.t0 42.3701
R87 Vp.n0 Vp.t3 39.1493
R88 Vp.n0 Vp.t2 38.876
R89 Vp Vp.n1 0.158324
R90 Vp Vp.n0 0.0370149
R91 GND.n31 GND.n6 109292
R92 GND.n34 GND.n31 50408.7
R93 GND.n21 GND.n10 37700.1
R94 GND.n90 GND.n89 15516.7
R95 GND.n88 GND.n10 10787.1
R96 GND.n79 GND.n70 8592.68
R97 GND.n73 GND.n70 8592.68
R98 GND.n79 GND.n71 8592.68
R99 GND.n73 GND.n71 8592.68
R100 GND.n61 GND.n22 8592.68
R101 GND.n57 GND.n22 8592.68
R102 GND.n61 GND.n23 8592.68
R103 GND.n57 GND.n23 8592.68
R104 GND.n42 GND.n30 6721.18
R105 GND.n42 GND.n35 6721.18
R106 GND.n38 GND.n30 6721.18
R107 GND.n96 GND.n7 6721.18
R108 GND.n91 GND.n7 6721.18
R109 GND.n96 GND.n8 6721.18
R110 GND.n91 GND.n8 6721.18
R111 GND.n33 GND.n29 5649.27
R112 GND.n47 GND.n29 5649.27
R113 GND.n47 GND.n28 5649.27
R114 GND.n33 GND.n28 5649.27
R115 GND.n100 GND.n4 4901.82
R116 GND.n100 GND.n5 4901.82
R117 GND.n101 GND.n4 4901.82
R118 GND.n101 GND.n5 4901.82
R119 GND.n82 GND.n12 4536.79
R120 GND.n86 GND.n12 4536.79
R121 GND.n82 GND.n13 4536.79
R122 GND.n86 GND.n13 4536.79
R123 GND.n64 GND.n17 4536.79
R124 GND.n68 GND.n17 4536.79
R125 GND.n64 GND.n18 4536.79
R126 GND.n68 GND.n18 4536.79
R127 GND.n89 GND.n9 3372.1
R128 GND.n10 GND.n9 2407.06
R129 GND.n44 GND.n30 2124.61
R130 GND.n31 GND.n9 1959.49
R131 GND.n44 GND.n34 1390.64
R132 GND.n88 GND.n87 1124.56
R133 GND.n44 GND.n43 844.298
R134 GND.n46 GND.n21 586.184
R135 GND.n58 GND.n56 558.307
R136 GND.n59 GND.n58 558.307
R137 GND.n74 GND.n72 558.307
R138 GND.n78 GND.n72 558.307
R139 GND.n45 GND.n44 554.826
R140 GND.n60 GND.n59 541.287
R141 GND.n78 GND.n77 537.958
R142 GND.n76 GND.n74 532.621
R143 GND.n98 GND.n97 509.024
R144 GND.n56 GND.n55 496.055
R145 GND.n41 GND.n40 436.707
R146 GND.n40 GND.n39 436.707
R147 GND.n93 GND.n92 436.707
R148 GND.n95 GND.n93 436.707
R149 GND.n95 GND.n94 434.397
R150 GND.n39 GND.n36 431.235
R151 GND.n92 GND.n1 428.851
R152 GND.n41 GND.n25 427.039
R153 GND.n63 GND.n21 368.741
R154 GND.n32 GND.n27 367.06
R155 GND.n32 GND.n26 367.06
R156 GND.n48 GND.n27 360.7
R157 GND.n49 GND.n26 359.651
R158 GND.n43 GND.t10 357.019
R159 GND.t4 GND.n45 357.019
R160 GND.t4 GND.n46 357.019
R161 GND.n38 GND.n37 343.635
R162 GND.n99 GND.n2 318.495
R163 GND.n99 GND.n3 318.495
R164 GND.n102 GND.n3 315.5
R165 GND.n103 GND.n2 313.651
R166 GND.n85 GND.n14 294.776
R167 GND.n85 GND.n84 294.776
R168 GND.n84 GND.n83 294.776
R169 GND.n67 GND.n19 294.776
R170 GND.n67 GND.n66 294.776
R171 GND.n66 GND.n65 294.776
R172 GND.n33 GND.n32 292.5
R173 GND.n34 GND.n33 292.5
R174 GND.n40 GND.n30 292.5
R175 GND.n48 GND.n47 292.5
R176 GND.n47 GND.t4 292.5
R177 GND.n36 GND.n35 292.5
R178 GND.n102 GND.n101 292.5
R179 GND.n101 GND.t0 292.5
R180 GND.n100 GND.n99 292.5
R181 GND.t0 GND.n100 292.5
R182 GND.n93 GND.n7 292.5
R183 GND.n7 GND.t11 292.5
R184 GND.n94 GND.n8 292.5
R185 GND.n8 GND.t11 292.5
R186 GND.n81 GND.n69 286.872
R187 GND.n37 GND.n35 265.971
R188 GND.n62 GND.t2 233.821
R189 GND.n80 GND.t6 233.821
R190 GND.t9 GND.n11 224.65
R191 GND.t8 GND.n16 216.792
R192 GND.n83 GND.n15 185.225
R193 GND.n65 GND.n20 177.683
R194 GND.t0 GND.n6 150.672
R195 GND.t0 GND.n98 150.672
R196 GND.n97 GND.t11 150.672
R197 GND.n90 GND.t11 150.672
R198 GND.n89 GND.n88 121.823
R199 GND.n20 GND.n19 100.507
R200 GND.n15 GND.n14 83.9534
R201 GND.n69 GND.n16 82.5251
R202 GND.n87 GND.n11 74.6656
R203 GND.n59 GND.n23 73.1255
R204 GND.n23 GND.t2 73.1255
R205 GND.n56 GND.n22 73.1255
R206 GND.n22 GND.t2 73.1255
R207 GND.n77 GND.n71 73.1255
R208 GND.n71 GND.t6 73.1255
R209 GND.n72 GND.n70 73.1255
R210 GND.n70 GND.t6 73.1255
R211 GND.n68 GND.n67 73.1255
R212 GND.n69 GND.n68 73.1255
R213 GND.n65 GND.n64 73.1255
R214 GND.n64 GND.n63 73.1255
R215 GND.n86 GND.n85 73.1255
R216 GND.n87 GND.n86 73.1255
R217 GND.n83 GND.n82 73.1255
R218 GND.n82 GND.n81 73.1255
R219 GND.n81 GND.n80 56.3268
R220 GND.n66 GND.n18 53.1823
R221 GND.t8 GND.n18 53.1823
R222 GND.n19 GND.n17 53.1823
R223 GND.t8 GND.n17 53.1823
R224 GND.n84 GND.n13 53.1823
R225 GND.t9 GND.n13 53.1823
R226 GND.n14 GND.n12 53.1823
R227 GND.t9 GND.n12 53.1823
R228 GND.n63 GND.n62 48.4673
R229 GND.n50 GND.t5 43.0348
R230 GND.n104 GND.t1 42.7363
R231 GND.n52 GND.t3 41.5589
R232 GND.n75 GND.t7 41.4501
R233 GND.n5 GND.n3 30.79
R234 GND.n98 GND.n5 30.79
R235 GND.n4 GND.n2 30.79
R236 GND.n6 GND.n4 30.79
R237 GND.n29 GND.n27 25.4353
R238 GND.n46 GND.n29 25.4353
R239 GND.n28 GND.n26 25.4353
R240 GND.n45 GND.n28 25.4353
R241 GND.n42 GND.n41 20.8934
R242 GND.n43 GND.n42 20.8934
R243 GND.n39 GND.n38 20.8934
R244 GND.n92 GND.n91 20.8934
R245 GND.n91 GND.n90 20.8934
R246 GND.n96 GND.n95 20.8934
R247 GND.n97 GND.n96 20.8934
R248 GND.n58 GND.n57 18.8715
R249 GND.n57 GND.n16 18.8715
R250 GND.n61 GND.n60 18.8715
R251 GND.n62 GND.n61 18.8715
R252 GND.n74 GND.n73 18.8715
R253 GND.n73 GND.n11 18.8715
R254 GND.n79 GND.n78 18.8715
R255 GND.n80 GND.n79 18.8715
R256 GND.t2 GND.t8 17.0294
R257 GND.n37 GND.t10 14.9557
R258 GND.n24 GND.n15 14.5995
R259 GND.n24 GND.n20 13.9046
R260 GND.n60 GND.n55 9.73383
R261 GND.n51 GND.n25 9.43581
R262 GND.n105 GND.n1 9.35362
R263 GND.n104 GND.n103 9.3005
R264 GND.n50 GND.n49 9.3005
R265 GND.t6 GND.t9 9.1699
R266 GND.n106 GND.n0 4.31023
R267 GND.n94 GND.n1 3.49141
R268 GND.n55 GND.n54 3.45562
R269 GND.n106 GND.n105 3.23962
R270 GND.n76 GND.n75 3.1005
R271 GND.n53 GND.n51 2.79925
R272 GND.n36 GND.n25 1.82907
R273 GND.n77 GND.n76 1.4405
R274 GND.n54 GND.n53 1.37696
R275 GND.n103 GND.n102 1.16414
R276 GND.n54 GND.n24 1.03107
R277 GND.n49 GND.n48 0.457643
R278 GND.n52 GND.n0 0.421374
R279 GND.n105 GND.n104 0.345988
R280 GND.n53 GND.n52 0.207089
R281 GND.n51 GND.n50 0.191582
R282 GND GND.n106 0.155057
R283 GND.n75 GND.n0 0.114923
R284 G.n0 G.t2 710.75
R285 G.n0 G.t3 710.722
R286 G.n0 G.t1 33.5848
R287 G.n0 G.t0 25.8008
R288 D10.n8 D10.n2 6324.71
R289 D10.n6 D10.n5 6324.71
R290 D10.n5 D10.n4 714.823
R291 D10.n8 D10.n7 714.823
R292 D10.n9 D10.n1 674.635
R293 D10.n3 D10.n1 674.635
R294 D10.n3 D10.n0 653.207
R295 D10.n10 D10.n9 609.367
R296 D10 D10.t1 23.3757
R297 D10.n10 D10.n0 12.6321
R298 D10.n9 D10.n8 10.8829
R299 D10.n5 D10.n3 10.8829
R300 D10 D10.t2 9.05168
R301 D10.n6 D10.n1 5.78175
R302 D10.n2 D10.n0 5.78175
R303 D10.n4 D10.n2 5.12417
R304 D10.n7 D10.n6 5.12417
R305 D10 D10.n10 1.8605
R306 D10.n7 D10.t0 0.654401
R307 D10.n4 D10.t0 0.654401
R308 IN+.t0 IN+.t2 674.149
R309 IN+.t4 IN+.t0 674.149
R310 IN+.t1 IN+.t4 674.149
R311 IN+.t3 IN+.t1 674.149
R312 IN+ IN+.t3 337.546
R313 D1.n1 D1.t0 41.5662
R314 D1.n1 D1.t1 30.2625
R315 D1.n3 D1.t3 23.7094
R316 D1 D1.t5 23.6938
R317 D1.n2 D1.t4 23.6789
R318 D1.n0 D1.t6 23.6372
R319 D1 D1.t2 23.6236
R320 D1.n0 D1.n3 5.4541
R321 D1.n3 D1.n2 5.30625
R322 D1.n2 D1.n1 2.24937
R323 D1 D1.n0 1.6212
R324 w_1686_7818.n20 w_1686_7818.n17 20696.5
R325 w_1686_7818.n21 w_1686_7818.n17 20696.5
R326 w_1686_7818.n20 w_1686_7818.n18 20696.5
R327 w_1686_7818.n21 w_1686_7818.n18 20696.5
R328 w_1686_7818.n5 w_1686_7818.n2 20696.5
R329 w_1686_7818.n6 w_1686_7818.n2 20696.5
R330 w_1686_7818.n5 w_1686_7818.n3 20696.5
R331 w_1686_7818.n6 w_1686_7818.n3 20696.5
R332 w_1686_7818.t19 w_1686_7818.t15 3588.18
R333 w_1686_7818.t11 w_1686_7818.t19 3588.18
R334 w_1686_7818.t17 w_1686_7818.t11 3588.18
R335 w_1686_7818.t13 w_1686_7818.t17 3588.18
R336 w_1686_7818.t5 w_1686_7818.t3 3588.18
R337 w_1686_7818.t7 w_1686_7818.t5 3588.18
R338 w_1686_7818.t9 w_1686_7818.t7 3588.18
R339 w_1686_7818.t1 w_1686_7818.t9 3588.18
R340 w_1686_7818.n22 w_1686_7818.n16 2207.62
R341 w_1686_7818.n19 w_1686_7818.n16 2207.62
R342 w_1686_7818.n19 w_1686_7818.n15 2207.62
R343 w_1686_7818.n7 w_1686_7818.n1 2207.62
R344 w_1686_7818.n4 w_1686_7818.n1 2207.62
R345 w_1686_7818.n4 w_1686_7818.n0 2207.62
R346 w_1686_7818.t15 w_1686_7818.n20 1908.11
R347 w_1686_7818.n21 w_1686_7818.t13 1908.11
R348 w_1686_7818.t3 w_1686_7818.n5 1908.11
R349 w_1686_7818.n6 w_1686_7818.t1 1908.11
R350 w_1686_7818.n23 w_1686_7818.n15 1617.86
R351 w_1686_7818.n8 w_1686_7818.n0 1565.89
R352 w_1686_7818.n23 w_1686_7818.n22 463.599
R353 w_1686_7818.n8 w_1686_7818.n7 429.7
R354 w_1686_7818.n25 w_1686_7818.t0 48.1635
R355 w_1686_7818.n22 w_1686_7818.n21 37.0005
R356 w_1686_7818.n20 w_1686_7818.n19 37.0005
R357 w_1686_7818.n7 w_1686_7818.n6 37.0005
R358 w_1686_7818.n5 w_1686_7818.n4 37.0005
R359 w_1686_7818.n9 w_1686_7818.t2 23.3782
R360 w_1686_7818.n24 w_1686_7818.t14 23.375
R361 w_1686_7818.n27 w_1686_7818.t12 23.3739
R362 w_1686_7818.n26 w_1686_7818.t18 23.3739
R363 w_1686_7818.n14 w_1686_7818.t16 23.3739
R364 w_1686_7818.n13 w_1686_7818.t4 23.3739
R365 w_1686_7818.n12 w_1686_7818.t6 23.3739
R366 w_1686_7818.n11 w_1686_7818.t8 23.3739
R367 w_1686_7818.n10 w_1686_7818.t10 23.3739
R368 w_1686_7818.t20 w_1686_7818.n28 23.3739
R369 w_1686_7818.n14 w_1686_7818.n13 1.71886
R370 w_1686_7818.n18 w_1686_7818.n16 1.12855
R371 w_1686_7818.t11 w_1686_7818.n18 1.12855
R372 w_1686_7818.n17 w_1686_7818.n15 1.12855
R373 w_1686_7818.t11 w_1686_7818.n17 1.12855
R374 w_1686_7818.n3 w_1686_7818.n1 1.12855
R375 w_1686_7818.t7 w_1686_7818.n3 1.12855
R376 w_1686_7818.n2 w_1686_7818.n0 1.12855
R377 w_1686_7818.t7 w_1686_7818.n2 1.12855
R378 w_1686_7818.n24 w_1686_7818.n23 1.03383
R379 w_1686_7818.n28 w_1686_7818.n14 0.532923
R380 w_1686_7818.n28 w_1686_7818.n27 0.531703
R381 w_1686_7818.n27 w_1686_7818.n26 0.528832
R382 w_1686_7818.n26 w_1686_7818.n25 0.423635
R383 w_1686_7818.n9 w_1686_7818.n8 0.423227
R384 w_1686_7818.n11 w_1686_7818.n10 0.422018
R385 w_1686_7818.n12 w_1686_7818.n11 0.415018
R386 w_1686_7818.n13 w_1686_7818.n12 0.414479
R387 w_1686_7818.n10 w_1686_7818.n9 0.403693
R388 w_1686_7818.n25 w_1686_7818.n24 0.243687
R389 Vc.t3 Vc.t4 126.523
R390 Vc.n1 Vc.t6 75.1209
R391 Vc.n4 Vc.t5 75.0448
R392 Vc.n7 Vc.t3 63.4118
R393 Vc.n0 Vc.t1 43.3772
R394 Vc.n0 Vc.t0 42.3701
R395 Vc.n2 Vc.t7 11.7318
R396 Vc.n3 Vc.t2 11.7318
R397 Vc.n7 Vc.n6 2.56155
R398 Vc.n5 Vc.n3 0.549556
R399 Vc Vc.n7 0.26415
R400 Vc.n1 Vc 0.23112
R401 Vc.n2 Vc 0.104667
R402 Vc.n4 Vc 0.0896473
R403 Vc.n4 Vc 0.0803267
R404 Vc.n6 Vc.n1 0.0697829
R405 Vc.n5 Vc.n4 0.0697829
R406 Vc.n6 Vc.n5 0.00340698
R407 Vc Vc.n0 0.0027007
R408 Vc.n3 Vc.n2 0.00216667
R409 IN-.t2 IN-.t1 674.284
R410 IN-.t3 IN-.t2 674.284
R411 IN-.t4 IN-.t3 674.284
R412 IN-.t0 IN-.t4 674.284
R413 IN- IN-.t0 337.548
R414 D2.n5 D2.t6 41.5839
R415 D2.n5 D2.t5 30.2422
R416 D2.n0 D2.t0 23.3739
R417 D2.n4 D2.t1 23.3739
R418 D2.n3 D2.t2 23.3739
R419 D2.n2 D2.t3 23.3739
R420 D2.n1 D2.t4 23.3739
R421 D2.n6 D2 3.10954
R422 D2.n2 D2 2.84864
R423 D2.n6 D2.n5 2.26609
R424 D2.n3 D2 2.23241
R425 D2.n4 D2 1.61947
R426 D2.n7 D2 1.40345
R427 D2.n8 D2 1.05044
R428 D2.n0 D2 1.00214
R429 D2.n9 D2 0.699307
R430 D2 D2.n1 0.425883
R431 D2.n1 D2 0.398526
R432 D2.n2 D2.n6 0.35686
R433 D2.n1 D2 0.34158
R434 D2.n1 D2.n0 0.233226
R435 D2.n9 D2.n4 0.229143
R436 D2.n8 D2.n3 0.229143
R437 D2.n7 D2.n2 0.229143
R438 D2.n0 D2.n9 0.218702
R439 D2.n3 D2.n7 0.217605
R440 D2.n4 D2.n8 0.214316
R441 D9.n9 D9.n8 6324.71
R442 D9.n6 D9.n4 6324.71
R443 D9.n4 D9.n3 714.823
R444 D9.n8 D9.n7 714.823
R445 D9.n5 D9.n2 674.635
R446 D9.n5 D9.n1 674.635
R447 D9.n0 D9.n2 637.811
R448 D9.n0 D9.n1 637.226
R449 D9 D9.t1 23.3739
R450 D9.n8 D9.n2 10.8829
R451 D9.n4 D9.n1 10.8829
R452 D9 D9.t2 9.05168
R453 D9.n6 D9.n5 5.78175
R454 D9.n0 D9.n9 5.78175
R455 D9.n9 D9.n3 5.12417
R456 D9.n7 D9.n6 5.12417
R457 D9 D9.n0 2.02907
R458 D9.n7 D9.t0 0.654401
R459 D9.t0 D9.n3 0.654401
R460 OUT.n0 OUT.t0 30.7611
R461 OUT.n0 OUT.t1 24.507
R462 OUT OUT.n0 4.84232
C0 D1 Vc 0.291331f
C1 D10 VDD 3.27648f
C2 a_3651_12640# VDD 0.998846f
C3 Vp D9 6.24e-20
C4 D2 OUT 0.797265f
C5 D9 Vc 2.2279f
C6 IN+ VDD 0.001874f
C7 Vp a_3651_12640# 0.454875f
C8 D1 IN+ 1.36571f
C9 D10 Vc 2.45204f
C10 D1 D2 1.22193f
C11 D1 VDD 0.006133f
C12 OUT Vc 2.67824f
C13 D9 IN+ 1.86e-19
C14 Vp VDD 4.52634f
C15 D9 VDD 3.27005f
C16 D10 OUT 0.97438f
C17 D1 Vp 0.004f
C18 D2 IN- 1.21532f
C19 D2 Vc 2.86656f
C20 VDD Vc 0.169798f
C21 D1 IN- 0.036349f
C22 IN- GND 4.018092f
C23 IN+ GND 4.048183f
C24 OUT GND 9.226859f
C25 VDD GND 54.74122f
C26 D2 GND 2.012658f
C27 D1 GND 12.38512f
C28 Vc GND 29.066322f
C29 a_3651_12640# GND 0.664555f
C30 Vp GND 6.420079f
C31 D10 GND 14.300781f
C32 D9 GND 14.618061f
C33 OUT.t1 GND 0.102957f
C34 OUT.t0 GND 0.02426f
C35 OUT.n0 GND 1.54873f
C36 D9.n0 GND 0.079161f
C37 D9.n1 GND 0.060212f
C38 D9.n2 GND 0.060236f
C39 D9.t0 GND 1.64637f
C40 D9.n4 GND 0.934717f
C41 D9.n5 GND 0.06131f
C42 D9.n6 GND 0.06131f
C43 D9.n8 GND 0.934717f
C44 D9.n9 GND 0.06131f
C45 D9.t1 GND 0.106336f
C46 D9.t2 GND 0.270761f
C47 D2.n0 GND 1.44819f
C48 D2.n1 GND 2.05847f
C49 D2.n2 GND 2.68057f
C50 D2.n3 GND 2.20807f
C51 D2.n4 GND 1.8259f
C52 D2.t5 GND 0.022985f
C53 D2.t6 GND 0.015218f
C54 D2.n5 GND 0.968435f
C55 D2.n6 GND 5.54069f
C56 D2.t3 GND 0.079315f
C57 D2.n7 GND 2.99625f
C58 D2.t2 GND 0.079315f
C59 D2.n8 GND 2.33106f
C60 D2.t1 GND 0.079315f
C61 D2.n9 GND 1.67023f
C62 D2.t0 GND 0.079315f
C63 D2.t4 GND 0.079315f
C64 IN-.t1 GND 0.439111f
C65 IN-.t2 GND 0.451193f
C66 IN-.t3 GND 0.451193f
C67 IN-.t4 GND 0.451193f
C68 IN-.t0 GND 0.357187f
C69 Vc.t1 GND 0.012338f
C70 Vc.t0 GND 0.007959f
C71 Vc.n0 GND 0.447696f
C72 Vc.t6 GND 0.200274f
C73 Vc.n1 GND 0.143319f
C74 Vc.t7 GND 0.745776f
C75 Vc.n2 GND 0.447261f
C76 Vc.t2 GND 0.745776f
C77 Vc.n3 GND 0.740185f
C78 Vc.t5 GND 0.200209f
C79 Vc.n4 GND 0.107687f
C80 Vc.n5 GND 0.196275f
C81 Vc.n6 GND 0.855039f
C82 Vc.t4 GND 2.62406f
C83 Vc.t3 GND 2.28572f
C84 Vc.n7 GND 2.27701f
C85 w_1686_7818.t2 GND 0.080909f
C86 w_1686_7818.n0 GND 0.129892f
C87 w_1686_7818.n1 GND 0.15149f
C88 w_1686_7818.n2 GND 0.15149f
C89 w_1686_7818.n3 GND 0.15149f
C90 w_1686_7818.n4 GND 0.152301f
C91 w_1686_7818.n5 GND 0.432773f
C92 w_1686_7818.t3 GND 0.77051f
C93 w_1686_7818.t5 GND 1.00556f
C94 w_1686_7818.t7 GND 1.00556f
C95 w_1686_7818.t9 GND 1.00556f
C96 w_1686_7818.t1 GND 0.77051f
C97 w_1686_7818.n6 GND 0.432773f
C98 w_1686_7818.n7 GND 0.092818f
C99 w_1686_7818.n8 GND 0.134135f
C100 w_1686_7818.n9 GND 1.17477f
C101 w_1686_7818.t10 GND 0.080807f
C102 w_1686_7818.n10 GND 1.2979f
C103 w_1686_7818.t8 GND 0.080807f
C104 w_1686_7818.n11 GND 1.3033f
C105 w_1686_7818.t6 GND 0.080807f
C106 w_1686_7818.n12 GND 1.30546f
C107 w_1686_7818.t4 GND 0.080807f
C108 w_1686_7818.n13 GND 2.02106f
C109 w_1686_7818.t16 GND 0.080807f
C110 w_1686_7818.n14 GND 1.67363f
C111 w_1686_7818.t14 GND 0.08083f
C112 w_1686_7818.n15 GND 0.13147f
C113 w_1686_7818.n16 GND 0.15149f
C114 w_1686_7818.n17 GND 0.15149f
C115 w_1686_7818.n18 GND 0.15149f
C116 w_1686_7818.n19 GND 0.152301f
C117 w_1686_7818.n20 GND 0.432773f
C118 w_1686_7818.t15 GND 0.77051f
C119 w_1686_7818.t19 GND 1.00556f
C120 w_1686_7818.t11 GND 1.00556f
C121 w_1686_7818.t17 GND 1.00556f
C122 w_1686_7818.t13 GND 0.77051f
C123 w_1686_7818.n21 GND 0.432773f
C124 w_1686_7818.n22 GND 0.093207f
C125 w_1686_7818.n23 GND 0.097953f
C126 w_1686_7818.n24 GND 0.839418f
C127 w_1686_7818.t0 GND 0.040499f
C128 w_1686_7818.n25 GND 0.487406f
C129 w_1686_7818.t18 GND 0.080807f
C130 w_1686_7818.n26 GND 0.934809f
C131 w_1686_7818.t12 GND 0.080807f
C132 w_1686_7818.n27 GND 1.08745f
C133 w_1686_7818.n28 GND 1.08658f
C134 w_1686_7818.t20 GND 0.080807f
C135 D1.n0 GND 1.47738f
C136 D1.t5 GND 0.107059f
C137 D1.t1 GND 0.030643f
C138 D1.t0 GND 0.020238f
C139 D1.n1 GND 0.856564f
C140 D1.t4 GND 0.107099f
C141 D1.n2 GND 2.34917f
C142 D1.t3 GND 0.107023f
C143 D1.n3 GND 1.23314f
C144 D1.t6 GND 0.106912f
C145 D1.t2 GND 0.106767f
C146 IN+.t2 GND 0.43765f
C147 IN+.t0 GND 0.453636f
C148 IN+.t4 GND 0.453636f
C149 IN+.t1 GND 0.453766f
C150 IN+.t3 GND 0.35688f
C151 D10.t1 GND 0.093784f
C152 D10.t2 GND 0.238709f
C153 D10.n0 GND 0.034136f
C154 D10.n1 GND 0.054052f
C155 D10.n2 GND 0.054052f
C156 D10.t0 GND 1.45148f
C157 D10.n3 GND 0.053574f
C158 D10.n5 GND 0.824068f
C159 D10.n6 GND 0.054052f
C160 D10.n8 GND 0.824068f
C161 D10.n9 GND 0.051978f
C162 D10.n10 GND 0.036261f
C163 G.n0 GND 6.22074f
C164 G.t3 GND 0.938364f
C165 G.t2 GND 0.938378f
C166 G.t1 GND 0.107955f
C167 G.t0 GND 0.194568f
C168 Vp.t3 GND 0.921868f
C169 Vp.t2 GND 0.914498f
C170 Vp.n0 GND 2.04727f
C171 Vp.t1 GND 0.013112f
C172 Vp.t0 GND 0.009746f
C173 Vp.n1 GND 0.472122f
C174 VDD.t8 GND 0.00557f
C175 VDD.n0 GND 0.046354f
C176 VDD.n1 GND 0.051068f
C177 VDD.n2 GND 0.051068f
C178 VDD.t5 GND 0.82732f
C179 VDD.n3 GND 0.051567f
C180 VDD.n5 GND 0.474058f
C181 VDD.n6 GND 0.051068f
C182 VDD.n8 GND 0.474058f
C183 VDD.n9 GND 0.030081f
C184 VDD.n10 GND 0.029088f
C185 VDD.n11 GND 0.032966f
C186 VDD.n12 GND 0.051567f
C187 VDD.n13 GND 0.474058f
C188 VDD.n14 GND 0.474058f
C189 VDD.n15 GND 0.051068f
C190 VDD.n16 GND 0.051068f
C191 VDD.t2 GND 0.82732f
C192 VDD.n19 GND 0.051068f
C193 VDD.n20 GND 0.042852f
C194 VDD.n21 GND 0.035361f
C195 VDD.t7 GND 0.012483f
C196 VDD.n22 GND 0.936968f
C197 VDD.t3 GND 0.138159f
C198 VDD.n23 GND 1.46353f
C199 VDD.t6 GND 0.138159f
C200 VDD.n24 GND 1.47437f
C201 VDD.n25 GND 0.358011f
C202 VDD.n26 GND 0.021787f
C203 VDD.n27 GND 0.022148f
C204 VDD.n29 GND 0.022693f
C205 VDD.n30 GND 0.022711f
C206 VDD.n31 GND 0.290376f
C207 VDD.t4 GND 0.4857f
C208 VDD.n33 GND 0.022693f
C209 VDD.n34 GND 0.290376f
C210 VDD.n35 GND 0.015469f
C211 VDD.n36 GND 0.063987f
C212 VDD.n37 GND 0.021735f
C213 VDD.n38 GND 0.022169f
C214 VDD.n40 GND 0.022693f
C215 VDD.n41 GND 0.022711f
C216 VDD.n42 GND 0.290376f
C217 VDD.t0 GND 0.4857f
C218 VDD.n44 GND 0.022693f
C219 VDD.n45 GND 0.290376f
C220 VDD.n46 GND 0.015429f
C221 VDD.n47 GND 0.020559f
C222 VDD.n48 GND 0.773085f
C223 VDD.n49 GND 0.321128f
C224 VDD.t1 GND 0.027194f
C225 VDD.n50 GND 0.419685f
C226 VDD.n51 GND 0.550246f
.ends

