magic
tech sky130A
magscale 1 2
timestamp 1740999383
<< viali >>
rect 6074 14470 6276 14526
rect 16580 14434 16862 14520
rect 4794 13728 4874 14040
rect 8462 13378 8818 13454
rect 14406 13408 14762 13484
rect 1494 12498 1572 12542
rect 2306 12520 2384 12564
rect 18148 12446 18238 12502
rect 19014 12384 19104 12440
rect 4782 12014 4862 12326
rect 2602 10704 3222 10778
rect 15634 9400 15736 9502
rect 17022 9412 17116 9476
rect 2548 8318 3324 8442
rect 17126 7118 17222 7404
rect 15330 5990 15536 6070
<< metal1 >>
rect 18914 15120 19252 15122
rect 384 15118 3816 15120
rect 4502 15118 19352 15120
rect 384 14714 19352 15118
rect 1438 14270 1682 14714
rect 3782 14380 4532 14714
rect 5210 14376 5674 14714
rect 6022 14526 6320 14714
rect 6022 14470 6074 14526
rect 6276 14470 6320 14526
rect 6022 14462 6320 14470
rect 1506 14098 1568 14270
rect 2692 14054 3596 14214
rect 5206 14170 5674 14376
rect 7078 14374 10132 14714
rect 2692 13760 3594 14054
rect 4826 14052 5674 14170
rect 1854 13754 3594 13760
rect 4788 14040 5674 14052
rect 1854 13482 3596 13754
rect 4788 13728 4794 14040
rect 4874 13728 5674 14040
rect 4788 13716 5674 13728
rect 4826 13654 5674 13716
rect 1854 12956 2064 13482
rect 2692 13480 3596 13482
rect 2692 13478 3594 13480
rect 1526 12742 2064 12956
rect 1526 12730 2058 12742
rect 2230 12564 2452 12996
rect 1418 12542 1658 12550
rect 1418 12498 1494 12542
rect 1572 12498 1658 12542
rect 1418 12418 1658 12498
rect 2230 12520 2306 12564
rect 2384 12520 2452 12564
rect 2230 12468 2452 12520
rect 2692 12532 3122 13478
rect 3782 12678 4530 13316
rect 2230 12418 2450 12468
rect 996 12054 2450 12418
rect 996 11276 1426 12054
rect 2692 11802 3586 12532
rect 5206 12430 5674 13654
rect 7948 13454 9292 14106
rect 11212 14098 12030 14378
rect 13054 14346 16108 14714
rect 16532 14520 16908 14714
rect 16532 14434 16580 14520
rect 16862 14434 16908 14520
rect 16532 14426 16908 14434
rect 18950 14314 19260 14714
rect 11446 13508 11754 14098
rect 7948 13378 8462 13454
rect 8818 13378 9292 13454
rect 7948 13304 9292 13378
rect 11378 13284 11388 13508
rect 11826 13284 11836 13508
rect 13966 13484 15314 14088
rect 18186 13956 18760 13962
rect 13966 13408 14406 13484
rect 14762 13408 15314 13484
rect 13966 13328 15314 13408
rect 16708 13718 16882 13720
rect 17498 13718 18760 13956
rect 16708 13708 18760 13718
rect 16708 13410 17848 13708
rect 18186 13678 18760 13708
rect 16708 13188 16998 13410
rect 17404 13404 17848 13410
rect 9674 12494 13574 13096
rect 4806 12338 5674 12430
rect 15694 12414 17002 13188
rect 17404 12538 17666 13404
rect 16302 12412 17002 12414
rect 4776 12326 5674 12338
rect 4776 12014 4782 12326
rect 4862 12014 5674 12326
rect 17374 12290 17384 12538
rect 17684 12290 17694 12538
rect 18154 12514 18234 12966
rect 18538 12892 18760 13678
rect 18538 12604 19072 12892
rect 18096 12502 18308 12514
rect 18096 12446 18148 12502
rect 18238 12446 18308 12502
rect 18096 12324 18308 12446
rect 18970 12440 19166 12468
rect 18970 12384 19014 12440
rect 19104 12384 19166 12440
rect 18970 12324 19166 12384
rect 7988 12206 7998 12278
rect 9352 12206 9362 12278
rect 4776 12002 5674 12014
rect 4806 11904 5674 12002
rect 14148 12038 15558 12282
rect 18096 12256 19166 12324
rect 18096 12176 19168 12256
rect 14148 11844 16950 12038
rect 18098 12002 19168 12176
rect 2692 11796 3008 11802
rect 14148 11760 16952 11844
rect 3736 11378 4530 11632
rect 996 11132 1100 11276
rect 1308 11132 1426 11276
rect 996 11130 1426 11132
rect 2168 11376 6488 11378
rect 10998 11376 14180 11378
rect 2168 11044 14180 11376
rect 2172 10778 3636 11044
rect 392 10608 1618 10718
rect 2172 10704 2602 10778
rect 3222 10704 3636 10778
rect 2172 10628 3636 10704
rect 4374 10622 5838 11044
rect 6280 11042 14180 11044
rect 6616 10624 8080 11042
rect 8868 10624 10332 11042
rect 10998 11040 14180 11042
rect 16658 11110 16952 11760
rect 17810 11110 18276 11118
rect 11130 10622 12590 11040
rect 392 10404 1840 10608
rect 3944 10444 4058 10578
rect 6184 10448 6298 10582
rect 8422 10450 8536 10584
rect 10658 10450 10772 10584
rect 392 10292 1618 10404
rect 2200 10344 2210 10398
rect 3518 10344 3528 10398
rect 4510 10340 4520 10394
rect 5750 10340 5760 10394
rect 6710 10336 6720 10388
rect 7996 10336 8006 10388
rect 9004 10338 9014 10394
rect 10144 10338 10154 10394
rect 11186 10334 11196 10400
rect 12430 10334 12440 10400
rect 13782 9116 14174 11040
rect 16658 10684 18276 11110
rect 18466 11070 18864 12002
rect 18456 10760 18466 11070
rect 18864 10760 18874 11070
rect 15932 10120 15942 10382
rect 16284 10120 16294 10382
rect 15622 9502 15748 9508
rect 15622 9492 15634 9502
rect 15736 9492 15748 9502
rect 15622 9398 15632 9492
rect 15740 9398 15750 9492
rect 15622 9394 15748 9398
rect 15284 9300 15294 9366
rect 15594 9300 15604 9366
rect 15968 9218 16254 10120
rect 16658 9330 16952 10684
rect 17810 10012 18276 10684
rect 17810 9596 19722 10012
rect 17010 9480 17128 9482
rect 17008 9398 17018 9480
rect 17124 9398 17134 9480
rect 17820 9450 19722 9596
rect 2182 8660 14182 9116
rect 15778 8960 16402 9218
rect 2184 8442 3648 8660
rect 400 8216 1626 8334
rect 2184 8318 2548 8442
rect 3324 8318 3648 8442
rect 2184 8240 3648 8318
rect 4358 8238 5822 8660
rect 6636 8238 8100 8660
rect 8862 8238 10326 8660
rect 11084 8240 12548 8660
rect 14494 8428 14504 8638
rect 14744 8622 14754 8638
rect 15322 8622 15562 8886
rect 14744 8450 15562 8622
rect 14744 8428 14754 8450
rect 400 8016 1832 8216
rect 15322 8200 15562 8450
rect 3950 8068 4058 8168
rect 6190 8068 6298 8168
rect 8420 8074 8528 8174
rect 10658 8062 10766 8162
rect 400 7908 1626 8016
rect 2172 7668 3628 8000
rect 4348 7668 5830 7994
rect 6626 7668 8082 7988
rect 8862 7668 10318 7996
rect 11110 7668 12566 7992
rect 15962 7944 16248 8960
rect 16678 8640 16918 8890
rect 16666 8490 16676 8640
rect 16918 8490 16928 8640
rect 16678 8230 16904 8490
rect 2172 7660 14176 7668
rect 2172 7466 13876 7660
rect 996 7132 1076 7328
rect 1302 7132 1440 7328
rect 2176 7212 13876 7466
rect 13866 7198 13876 7212
rect 14514 7198 14524 7660
rect 996 5792 1440 7132
rect 15714 6426 16566 7944
rect 18456 7726 18466 8086
rect 18864 7726 18874 8086
rect 17120 7404 17228 7416
rect 17120 7118 17126 7404
rect 17222 7400 17228 7404
rect 17120 7112 17130 7118
rect 17232 7112 17242 7400
rect 17120 7106 17228 7112
rect 17356 6456 17366 6622
rect 17554 6620 17564 6622
rect 17554 6456 17596 6620
rect 15308 6070 15568 6154
rect 15308 5990 15330 6070
rect 15536 5990 15568 6070
rect 15308 5792 15568 5990
rect 16666 5792 16944 6186
rect 17356 5792 17596 6456
rect 18466 5798 18864 7726
rect 18466 5792 19366 5798
rect 404 5390 19366 5792
rect 404 5386 18602 5390
rect 996 5384 1440 5386
<< via1 >>
rect 11388 13284 11826 13508
rect 17384 12290 17684 12538
rect 7998 12206 9352 12278
rect 1100 11132 1308 11276
rect 2210 10344 3518 10398
rect 4520 10340 5750 10394
rect 6720 10336 7996 10388
rect 9014 10338 10144 10394
rect 11196 10334 12430 10400
rect 18466 10760 18864 11070
rect 15942 10120 16284 10382
rect 15632 9400 15634 9492
rect 15634 9400 15736 9492
rect 15736 9400 15740 9492
rect 15632 9398 15740 9400
rect 15294 9300 15594 9366
rect 17018 9476 17124 9480
rect 17018 9412 17022 9476
rect 17022 9412 17116 9476
rect 17116 9412 17124 9476
rect 17018 9398 17124 9412
rect 14504 8428 14744 8638
rect 16676 8490 16918 8640
rect 1076 7132 1302 7328
rect 13876 7198 14514 7660
rect 18466 7726 18864 8086
rect 17130 7118 17222 7400
rect 17222 7118 17232 7400
rect 17130 7112 17232 7118
rect 17366 6456 17554 6622
<< metal2 >>
rect 11388 13508 11826 13518
rect 11388 13274 11826 13284
rect 7998 12278 9352 12288
rect 7998 12196 9352 12206
rect 7998 11654 9342 12196
rect 7998 11652 10086 11654
rect 11444 11652 11790 13274
rect 17374 12538 17692 12548
rect 17374 12534 17384 12538
rect 17370 12290 17384 12534
rect 17684 12534 17692 12538
rect 17684 12290 17734 12534
rect 7998 11340 15598 11652
rect 7998 11338 10086 11340
rect 1100 11276 1308 11286
rect 1100 11130 1308 11132
rect 996 7328 1430 11130
rect 2210 10398 3518 10408
rect 2158 10344 2210 10380
rect 4520 10394 5750 10404
rect 3518 10344 3556 10380
rect 2158 9998 3556 10344
rect 4438 10340 4520 10384
rect 6720 10388 7996 10398
rect 5750 10340 5836 10384
rect 4438 9998 5836 10340
rect 6658 10336 6720 10386
rect 9014 10394 10144 10404
rect 7996 10336 8056 10386
rect 6658 10002 8056 10336
rect 8928 10338 9014 10384
rect 11196 10400 12430 10410
rect 10144 10338 10326 10384
rect 8928 10322 10326 10338
rect 11112 10334 11196 10392
rect 12430 10334 12518 10392
rect 8924 10016 10330 10322
rect 11112 10016 12518 10334
rect 8450 10002 13646 10016
rect 2156 9996 5892 9998
rect 6658 9996 13646 10002
rect 2156 9660 13646 9996
rect 8450 9654 13646 9660
rect 8924 9638 10330 9654
rect 13134 9608 13630 9654
rect 13128 8734 13632 9608
rect 15302 9376 15588 11340
rect 17370 10450 17734 12290
rect 18466 11070 18864 11080
rect 18864 10760 18874 11060
rect 18466 10750 18874 10760
rect 15940 10382 17734 10450
rect 15940 10120 15942 10382
rect 16284 10120 17734 10382
rect 15940 10056 17734 10120
rect 15622 9778 17482 9820
rect 15622 9570 17640 9778
rect 15622 9494 15764 9570
rect 15622 9492 15636 9494
rect 15734 9492 15764 9494
rect 15622 9448 15632 9492
rect 15740 9448 15764 9492
rect 16986 9480 17148 9570
rect 16986 9436 17018 9480
rect 15632 9388 15740 9398
rect 17124 9436 17148 9480
rect 17018 9388 17124 9398
rect 15294 9366 15594 9376
rect 15294 9290 15594 9300
rect 13128 8648 14740 8734
rect 13128 8638 14744 8648
rect 13128 8428 14504 8638
rect 16676 8640 16918 8650
rect 16676 8480 16918 8490
rect 13128 8418 14744 8428
rect 13128 8368 14740 8418
rect 996 7132 1076 7328
rect 1302 7132 1430 7328
rect 13876 7660 14514 7670
rect 17318 7494 17640 9570
rect 18476 9554 18874 10750
rect 18466 9262 18874 9554
rect 18466 8086 18864 9262
rect 18466 7716 18864 7726
rect 17138 7410 17644 7494
rect 13876 7188 14514 7198
rect 17130 7400 17644 7410
rect 17232 7112 17644 7400
rect 17130 7102 17644 7112
rect 17138 6966 17644 7102
rect 17318 6622 17640 6966
rect 17318 6456 17366 6622
rect 17554 6456 17640 6622
rect 17318 6436 17640 6456
<< via2 >>
rect 15636 9492 15734 9494
rect 15636 9398 15734 9492
rect 16676 8490 16918 8640
rect 13876 7198 14514 7660
<< metal3 >>
rect 13908 10342 14568 10352
rect 13908 10320 18020 10342
rect 13908 9782 18034 10320
rect 13908 9198 14568 9782
rect 15626 9494 15744 9499
rect 15626 9398 15636 9494
rect 15734 9398 15744 9494
rect 15626 9393 15744 9398
rect 13908 7665 14558 9198
rect 17546 8682 18034 9782
rect 16678 8645 18034 8682
rect 16666 8640 18034 8645
rect 16666 8490 16676 8640
rect 16918 8490 18034 8640
rect 16666 8485 18034 8490
rect 16678 8438 18034 8485
rect 13866 7660 14558 7665
rect 13866 7198 13876 7660
rect 14514 7198 14558 7660
rect 13866 7193 14558 7198
rect 13908 7188 14558 7193
use sky130_fd_pr__pfet_01v8_6HANBW  XM1
timestamp 1740997949
transform 0 1 7377 -1 0 10504
box -296 -5691 296 5691
use sky130_fd_pr__pfet_01v8_6HANBW  XM2
timestamp 1740997949
transform 0 1 7377 -1 0 8114
box -296 -5691 296 5691
use sky130_fd_pr__nfet_01v8_Q33MQV  XM3
timestamp 1740997949
transform 0 1 15442 -1 0 7176
box -1196 -410 1196 410
use sky130_fd_pr__nfet_01v8_Q33MQV  XM4
timestamp 1740997949
transform 0 1 16806 -1 0 7188
box -1196 -410 1196 410
use sky130_fd_pr__nfet_01v8_P3FTKA  XM5
timestamp 1740997949
transform 0 1 15428 -1 0 9100
box -396 -510 396 510
use sky130_fd_pr__nfet_01v8_P3FTKA  XM6
timestamp 1740997949
transform 0 1 16780 -1 0 9090
box -396 -510 396 510
use sky130_fd_pr__pfet_01v8_TKMKND  XM7
timestamp 1740997949
transform 0 1 8639 -1 0 12780
box -696 -1219 696 1219
use sky130_fd_pr__pfet_01v8_TKMKND  XM8
timestamp 1740997949
transform 0 1 14659 -1 0 12798
box -696 -1219 696 1219
use sky130_fd_pr__pfet_01v8_2C2MAW  XM9
timestamp 1740997949
transform 0 1 8613 -1 0 14248
box -296 -2769 296 2769
use sky130_fd_pr__pfet_01v8_2C2MAW  XM10
timestamp 1740997949
transform 0 1 14647 -1 0 14222
box -296 -2769 296 2769
use sky130_fd_pr__pfet_01v8_SKC8VM  XM11
timestamp 1740997949
transform 0 1 4151 -1 0 12140
box -696 -719 696 719
use sky130_fd_pr__pfet_01v8_SKC8VM  XM12
timestamp 1740997949
transform 0 1 4167 -1 0 13848
box -696 -719 696 719
use sky130_fd_pr__res_xhigh_po_0p35_8HWFQE  XR1
timestamp 1740997949
transform 1 0 18191 0 1 13323
box -201 -897 201 897
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR2
timestamp 1740997949
transform 1 0 1545 0 1 13552
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_YTZ25J  XR3
timestamp 1740997949
transform 1 0 2341 0 1 13256
box -201 -768 201 768
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR5
timestamp 1740997949
transform 1 0 19067 0 1 13438
box -201 -1082 201 1082
<< labels >>
flabel metal1 472 8016 672 8216 0 FreeSans 256 0 0 0 IN-
port 3 nsew
flabel metal1 494 5486 694 5686 0 FreeSans 256 0 0 0 GND
port 1 nsew
flabel metal1 482 14838 682 15038 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 480 10406 680 10606 0 FreeSans 256 0 0 0 IN+
port 2 nsew
flabel metal1 19344 9624 19544 9824 0 FreeSans 256 0 0 0 OUT
port 4 nsew
rlabel metal1 2692 13478 3594 14214 1 Vp
rlabel metal1 18186 13678 18760 13962 1 Vc
rlabel metal1 11446 13508 11754 14378 1 G
rlabel metal2 2158 9660 3556 10344 1 D1
rlabel metal1 2176 7212 13876 7668 1 D2
rlabel metal1 7948 13454 9292 14106 1 D9
rlabel metal1 13966 13484 15314 14088 1 D10
rlabel metal1 15778 8960 16402 9218 1 Vc
rlabel metal1 15714 6426 16566 7944 1 Vc
rlabel space 3736 11044 4530 11634 1 S
<< end >>
