magic
tech sky130A
magscale 1 2
timestamp 1741188478
<< nwell >>
rect -296 -5691 296 5691
<< pmos >>
rect -100 3472 100 5472
rect -100 1236 100 3236
rect -100 -1000 100 1000
rect -100 -3236 100 -1236
rect -100 -5472 100 -3472
<< pdiff >>
rect -158 5460 -100 5472
rect -158 3484 -146 5460
rect -112 3484 -100 5460
rect -158 3472 -100 3484
rect 100 5460 158 5472
rect 100 3484 112 5460
rect 146 3484 158 5460
rect 100 3472 158 3484
rect -158 3224 -100 3236
rect -158 1248 -146 3224
rect -112 1248 -100 3224
rect -158 1236 -100 1248
rect 100 3224 158 3236
rect 100 1248 112 3224
rect 146 1248 158 3224
rect 100 1236 158 1248
rect -158 988 -100 1000
rect -158 -988 -146 988
rect -112 -988 -100 988
rect -158 -1000 -100 -988
rect 100 988 158 1000
rect 100 -988 112 988
rect 146 -988 158 988
rect 100 -1000 158 -988
rect -158 -1248 -100 -1236
rect -158 -3224 -146 -1248
rect -112 -3224 -100 -1248
rect -158 -3236 -100 -3224
rect 100 -1248 158 -1236
rect 100 -3224 112 -1248
rect 146 -3224 158 -1248
rect 100 -3236 158 -3224
rect -158 -3484 -100 -3472
rect -158 -5460 -146 -3484
rect -112 -5460 -100 -3484
rect -158 -5472 -100 -5460
rect 100 -3484 158 -3472
rect 100 -5460 112 -3484
rect 146 -5460 158 -3484
rect 100 -5472 158 -5460
<< pdiffc >>
rect -146 3484 -112 5460
rect 112 3484 146 5460
rect -146 1248 -112 3224
rect 112 1248 146 3224
rect -146 -988 -112 988
rect 112 -988 146 988
rect -146 -3224 -112 -1248
rect 112 -3224 146 -1248
rect -146 -5460 -112 -3484
rect 112 -5460 146 -3484
<< nsubdiff >>
rect -260 5621 -164 5655
rect 164 5621 260 5655
rect -260 5559 -226 5621
rect 226 5559 260 5621
rect -260 -5621 -226 -5559
rect 226 -5621 260 -5559
rect -260 -5655 -164 -5621
rect 164 -5655 260 -5621
<< nsubdiffcont >>
rect -164 5621 164 5655
rect -260 -5559 -226 5559
rect 226 -5559 260 5559
rect -164 -5655 164 -5621
<< poly >>
rect -100 5553 100 5569
rect -100 5519 -84 5553
rect 84 5519 100 5553
rect -100 5472 100 5519
rect -100 3425 100 3472
rect -100 3391 -84 3425
rect 84 3391 100 3425
rect -100 3375 100 3391
rect -100 3317 100 3333
rect -100 3283 -84 3317
rect 84 3283 100 3317
rect -100 3236 100 3283
rect -100 1189 100 1236
rect -100 1155 -84 1189
rect 84 1155 100 1189
rect -100 1139 100 1155
rect -100 1081 100 1097
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -100 1000 100 1047
rect -100 -1047 100 -1000
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1097 100 -1081
rect -100 -1155 100 -1139
rect -100 -1189 -84 -1155
rect 84 -1189 100 -1155
rect -100 -1236 100 -1189
rect -100 -3283 100 -3236
rect -100 -3317 -84 -3283
rect 84 -3317 100 -3283
rect -100 -3333 100 -3317
rect -100 -3391 100 -3375
rect -100 -3425 -84 -3391
rect 84 -3425 100 -3391
rect -100 -3472 100 -3425
rect -100 -5519 100 -5472
rect -100 -5553 -84 -5519
rect 84 -5553 100 -5519
rect -100 -5569 100 -5553
<< polycont >>
rect -84 5519 84 5553
rect -84 3391 84 3425
rect -84 3283 84 3317
rect -84 1155 84 1189
rect -84 1047 84 1081
rect -84 -1081 84 -1047
rect -84 -1189 84 -1155
rect -84 -3317 84 -3283
rect -84 -3425 84 -3391
rect -84 -5553 84 -5519
<< locali >>
rect -260 5621 -164 5655
rect 164 5621 260 5655
rect -260 5559 -226 5621
rect 226 5559 260 5621
rect -100 5519 -84 5553
rect 84 5519 100 5553
rect -146 5460 -112 5476
rect -146 3468 -112 3484
rect 112 5460 146 5476
rect 112 3468 146 3484
rect -100 3391 -84 3425
rect 84 3391 100 3425
rect -100 3283 -84 3317
rect 84 3283 100 3317
rect -146 3224 -112 3240
rect -146 1232 -112 1248
rect 112 3224 146 3240
rect 112 1232 146 1248
rect -100 1155 -84 1189
rect 84 1155 100 1189
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -146 988 -112 1004
rect -146 -1004 -112 -988
rect 112 988 146 1004
rect 112 -1004 146 -988
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1189 -84 -1155
rect 84 -1189 100 -1155
rect -146 -1248 -112 -1232
rect -146 -3240 -112 -3224
rect 112 -1248 146 -1232
rect 112 -3240 146 -3224
rect -100 -3317 -84 -3283
rect 84 -3317 100 -3283
rect -100 -3425 -84 -3391
rect 84 -3425 100 -3391
rect -146 -3484 -112 -3468
rect -146 -5476 -112 -5460
rect 112 -3484 146 -3468
rect 112 -5476 146 -5460
rect -100 -5553 -84 -5519
rect 84 -5553 100 -5519
rect -260 -5621 -226 -5559
rect 226 -5621 260 -5559
rect -260 -5655 -164 -5621
rect 164 -5655 260 -5621
<< viali >>
rect -84 5519 84 5553
rect -146 3484 -112 5460
rect 112 3484 146 5460
rect -84 3391 84 3425
rect -84 3283 84 3317
rect -146 1248 -112 3224
rect 112 1248 146 3224
rect -84 1155 84 1189
rect -84 1047 84 1081
rect -146 -988 -112 988
rect 112 -988 146 988
rect -84 -1081 84 -1047
rect -84 -1189 84 -1155
rect -146 -3224 -112 -1248
rect 112 -3224 146 -1248
rect -84 -3317 84 -3283
rect -84 -3425 84 -3391
rect -146 -5460 -112 -3484
rect 112 -5460 146 -3484
rect -84 -5553 84 -5519
<< metal1 >>
rect -96 5553 96 5559
rect -96 5519 -84 5553
rect 84 5519 96 5553
rect -96 5513 96 5519
rect -152 5460 -106 5472
rect -152 3484 -146 5460
rect -112 3484 -106 5460
rect -152 3472 -106 3484
rect 106 5460 152 5472
rect 106 3484 112 5460
rect 146 3484 152 5460
rect 106 3472 152 3484
rect -96 3425 96 3431
rect -96 3391 -84 3425
rect 84 3391 96 3425
rect -96 3385 96 3391
rect -96 3317 96 3323
rect -96 3283 -84 3317
rect 84 3283 96 3317
rect -96 3277 96 3283
rect -152 3224 -106 3236
rect -152 1248 -146 3224
rect -112 1248 -106 3224
rect -152 1236 -106 1248
rect 106 3224 152 3236
rect 106 1248 112 3224
rect 146 1248 152 3224
rect 106 1236 152 1248
rect -96 1189 96 1195
rect -96 1155 -84 1189
rect 84 1155 96 1189
rect -96 1149 96 1155
rect -96 1081 96 1087
rect -96 1047 -84 1081
rect 84 1047 96 1081
rect -96 1041 96 1047
rect -152 988 -106 1000
rect -152 -988 -146 988
rect -112 -988 -106 988
rect -152 -1000 -106 -988
rect 106 988 152 1000
rect 106 -988 112 988
rect 146 -988 152 988
rect 106 -1000 152 -988
rect -96 -1047 96 -1041
rect -96 -1081 -84 -1047
rect 84 -1081 96 -1047
rect -96 -1087 96 -1081
rect -96 -1155 96 -1149
rect -96 -1189 -84 -1155
rect 84 -1189 96 -1155
rect -96 -1195 96 -1189
rect -152 -1248 -106 -1236
rect -152 -3224 -146 -1248
rect -112 -3224 -106 -1248
rect -152 -3236 -106 -3224
rect 106 -1248 152 -1236
rect 106 -3224 112 -1248
rect 146 -3224 152 -1248
rect 106 -3236 152 -3224
rect -96 -3283 96 -3277
rect -96 -3317 -84 -3283
rect 84 -3317 96 -3283
rect -96 -3323 96 -3317
rect -96 -3391 96 -3385
rect -96 -3425 -84 -3391
rect 84 -3425 96 -3391
rect -96 -3431 96 -3425
rect -152 -3484 -106 -3472
rect -152 -5460 -146 -3484
rect -112 -5460 -106 -3484
rect -152 -5472 -106 -5460
rect 106 -3484 152 -3472
rect 106 -5460 112 -3484
rect 146 -5460 152 -3484
rect 106 -5472 152 -5460
rect -96 -5519 96 -5513
rect -96 -5553 -84 -5519
rect 84 -5553 96 -5519
rect -96 -5559 96 -5553
<< properties >>
string FIXED_BBOX -243 -5638 243 5638
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
