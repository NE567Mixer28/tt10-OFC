magic
tech sky130A
magscale 1 2
timestamp 1741188478
<< pwell >>
rect -201 -897 201 897
<< psubdiff >>
rect -165 827 -69 861
rect 69 827 165 861
rect -165 765 -131 827
rect 131 765 165 827
rect -165 -827 -131 -765
rect 131 -827 165 -765
rect -165 -861 -69 -827
rect 69 -861 165 -827
<< psubdiffcont >>
rect -69 827 69 861
rect -165 -765 -131 765
rect 131 -765 165 765
rect -69 -861 69 -827
<< xpolycontact >>
rect -35 299 35 731
rect -35 -731 35 -299
<< xpolyres >>
rect -35 -299 35 299
<< locali >>
rect -165 827 -69 861
rect 69 827 165 861
rect -165 765 -131 827
rect 131 765 165 827
rect -165 -827 -131 -765
rect 131 -827 165 -765
rect -165 -861 -69 -827
rect 69 -861 165 -827
<< viali >>
rect -19 316 19 713
rect -19 -713 19 -316
<< metal1 >>
rect -25 713 25 725
rect -25 316 -19 713
rect 19 316 25 713
rect -25 304 25 316
rect -25 -316 25 -304
rect -25 -713 -19 -316
rect 19 -713 25 -316
rect -25 -725 25 -713
<< properties >>
string FIXED_BBOX -148 -844 148 844
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 3.15 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 19.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
